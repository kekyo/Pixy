module Core(
	output SRAMCS0,
	output SRAMCS1,
	output PROMCS0,
	output PROMCS1
);

assign SRAMCS0 = 0;
assign SRAMCS1 = 0;
assign PROMCS0 = 0;
assign PROMCS1 = 0;

endmodule